LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INVERSORA IS
PORT(X: in std_logic;
	Y: out std_logic);
END INVERSORA;

ARCHITECTURE INVERSORA_ARCH OF INVERSORA IS
BEGIN
	Y <= not(X);

END INVERSORA_ARCH;